module tb_fifo;
    bit clk;
    bit ref_clk;